--==============================================================================
-- Project: Pixel Processing
-- Author : Kevin Hughes
-- Date   : Monday, December 17th, 2018
-- Module : lookup_table.vhd
-- Desc.  : Calculates the vertical Sobel output of a given matrix.
--==============================================================================
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--==============================================================================
-- LOOKUP_TABLE Entity Block
-- I_EDGE_VALUE : Combined edge detection magnitude squared
-- O_PIX_VALUE  : Combined edge detection magnitude
--==============================================================================
entity LOOKUP_TABLE is
port(
	I_EDGE_VALUE : in std_logic_vector(20 downto 0);
	O_PIX_VALUE  : out std_logic_vector(7 downto 0)
);end entity LOOKUP_TABLE;

--==============================================================================
-- LOOKUP_TABLE Architecture Block
--==============================================================================
architecture RTL of LOOKUP_TABLE is

signal INT_EDGE_VALUE : integer; 

begin

INT_EDGE_VALUE <= to_integer(unsigned(I_EDGE_VALUE));

O_PIX_VALUE <= 
"00000000" when INT_EDGE_VALUE <= 7 else 
"00000001" when INT_EDGE_VALUE >= 8 and INT_EDGE_VALUE <= 72 else 
"00000010" when INT_EDGE_VALUE >= 73 and INT_EDGE_VALUE <= 199 else 
"00000011" when INT_EDGE_VALUE >= 200 and INT_EDGE_VALUE <= 391 else 
"00000100" when INT_EDGE_VALUE >= 392 and INT_EDGE_VALUE <= 647 else 
"00000101" when INT_EDGE_VALUE >= 648 and INT_EDGE_VALUE <= 967 else 
"00000110" when INT_EDGE_VALUE >= 968 and INT_EDGE_VALUE <= 1351 else 
"00000111" when INT_EDGE_VALUE >= 1352 and INT_EDGE_VALUE <= 1799 else 
"00001000" when INT_EDGE_VALUE >= 1800 and INT_EDGE_VALUE <= 2311 else 
"00001001" when INT_EDGE_VALUE >= 2312 and INT_EDGE_VALUE <= 2887 else 
"00001010" when INT_EDGE_VALUE >= 2888 and INT_EDGE_VALUE <= 3527 else 
"00001011" when INT_EDGE_VALUE >= 3528 and INT_EDGE_VALUE <= 4231 else 
"00001100" when INT_EDGE_VALUE >= 4232 and INT_EDGE_VALUE <= 4999 else 
"00001101" when INT_EDGE_VALUE >= 5000 and INT_EDGE_VALUE <= 5831 else 
"00001110" when INT_EDGE_VALUE >= 5832 and INT_EDGE_VALUE <= 6728 else 
"00001111" when INT_EDGE_VALUE >= 6729 and INT_EDGE_VALUE <= 7687 else 
"00010000" when INT_EDGE_VALUE >= 7688 and INT_EDGE_VALUE <= 8712 else 
"00010001" when INT_EDGE_VALUE >= 8713 and INT_EDGE_VALUE <= 9799 else 
"00010010" when INT_EDGE_VALUE >= 9800 and INT_EDGE_VALUE <= 10951 else 
"00010011" when INT_EDGE_VALUE >= 10952 and INT_EDGE_VALUE <= 12168 else 
"00010100" when INT_EDGE_VALUE >= 12169 and INT_EDGE_VALUE <= 13448 else 
"00010101" when INT_EDGE_VALUE >= 13449 and INT_EDGE_VALUE <= 14792 else 
"00010110" when INT_EDGE_VALUE >= 14793 and INT_EDGE_VALUE <= 16199 else 
"00010111" when INT_EDGE_VALUE >= 16200 and INT_EDGE_VALUE <= 17672 else 
"00011000" when INT_EDGE_VALUE >= 17673 and INT_EDGE_VALUE <= 19207 else 
"00011001" when INT_EDGE_VALUE >= 19208 and INT_EDGE_VALUE <= 20808 else 
"00011010" when INT_EDGE_VALUE >= 20809 and INT_EDGE_VALUE <= 22472 else 
"00011011" when INT_EDGE_VALUE >= 22473 and INT_EDGE_VALUE <= 24199 else 
"00011100" when INT_EDGE_VALUE >= 24200 and INT_EDGE_VALUE <= 25992 else 
"00011101" when INT_EDGE_VALUE >= 25993 and INT_EDGE_VALUE <= 27847 else 
"00011110" when INT_EDGE_VALUE >= 27848 and INT_EDGE_VALUE <= 29768 else 
"00011111" when INT_EDGE_VALUE >= 29769 and INT_EDGE_VALUE <= 31752 else 
"00100000" when INT_EDGE_VALUE >= 31753 and INT_EDGE_VALUE <= 33799 else 
"00100001" when INT_EDGE_VALUE >= 33800 and INT_EDGE_VALUE <= 35911 else 
"00100010" when INT_EDGE_VALUE >= 35912 and INT_EDGE_VALUE <= 38087 else 
"00100011" when INT_EDGE_VALUE >= 38088 and INT_EDGE_VALUE <= 40327 else 
"00100100" when INT_EDGE_VALUE >= 40328 and INT_EDGE_VALUE <= 42631 else 
"00100101" when INT_EDGE_VALUE >= 42632 and INT_EDGE_VALUE <= 44999 else 
"00100110" when INT_EDGE_VALUE >= 45000 and INT_EDGE_VALUE <= 47431 else 
"00100111" when INT_EDGE_VALUE >= 47432 and INT_EDGE_VALUE <= 49927 else 
"00101000" when INT_EDGE_VALUE >= 49928 and INT_EDGE_VALUE <= 52487 else 
"00101001" when INT_EDGE_VALUE >= 52488 and INT_EDGE_VALUE <= 55112 else 
"00101010" when INT_EDGE_VALUE >= 55113 and INT_EDGE_VALUE <= 57799 else 
"00101011" when INT_EDGE_VALUE >= 57800 and INT_EDGE_VALUE <= 60551 else 
"00101100" when INT_EDGE_VALUE >= 60552 and INT_EDGE_VALUE <= 63367 else 
"00101101" when INT_EDGE_VALUE >= 63368 and INT_EDGE_VALUE <= 66248 else 
"00101110" when INT_EDGE_VALUE >= 66249 and INT_EDGE_VALUE <= 69191 else 
"00101111" when INT_EDGE_VALUE >= 69192 and INT_EDGE_VALUE <= 72199 else 
"00110000" when INT_EDGE_VALUE >= 72200 and INT_EDGE_VALUE <= 75271 else 
"00110001" when INT_EDGE_VALUE >= 75272 and INT_EDGE_VALUE <= 78408 else 
"00110010" when INT_EDGE_VALUE >= 78409 and INT_EDGE_VALUE <= 81608 else 
"00110011" when INT_EDGE_VALUE >= 81609 and INT_EDGE_VALUE <= 84871 else 
"00110100" when INT_EDGE_VALUE >= 84872 and INT_EDGE_VALUE <= 88199 else 
"00110101" when INT_EDGE_VALUE >= 88200 and INT_EDGE_VALUE <= 91591 else 
"00110110" when INT_EDGE_VALUE >= 91592 and INT_EDGE_VALUE <= 95047 else 
"00110111" when INT_EDGE_VALUE >= 95048 and INT_EDGE_VALUE <= 98568 else 
"00111000" when INT_EDGE_VALUE >= 98569 and INT_EDGE_VALUE <= 102151 else 
"00111001" when INT_EDGE_VALUE >= 102152 and INT_EDGE_VALUE <= 105799 else 
"00111010" when INT_EDGE_VALUE >= 105800 and INT_EDGE_VALUE <= 109511 else 
"00111011" when INT_EDGE_VALUE >= 109512 and INT_EDGE_VALUE <= 113288 else 
"00111100" when INT_EDGE_VALUE >= 113289 and INT_EDGE_VALUE <= 117127 else 
"00111101" when INT_EDGE_VALUE >= 117128 and INT_EDGE_VALUE <= 121031 else 
"00111110" when INT_EDGE_VALUE >= 121032 and INT_EDGE_VALUE <= 124999 else 
"00111111" when INT_EDGE_VALUE >= 125000 and INT_EDGE_VALUE <= 129031 else 
"01000000" when INT_EDGE_VALUE >= 129032 and INT_EDGE_VALUE <= 133127 else 
"01000001" when INT_EDGE_VALUE >= 133128 and INT_EDGE_VALUE <= 137287 else 
"01000010" when INT_EDGE_VALUE >= 137288 and INT_EDGE_VALUE <= 141511 else 
"01000011" when INT_EDGE_VALUE >= 141512 and INT_EDGE_VALUE <= 145799 else 
"01000100" when INT_EDGE_VALUE >= 145800 and INT_EDGE_VALUE <= 150151 else 
"01000101" when INT_EDGE_VALUE >= 150152 and INT_EDGE_VALUE <= 154567 else 
"01000110" when INT_EDGE_VALUE >= 154568 and INT_EDGE_VALUE <= 159048 else 
"01000111" when INT_EDGE_VALUE >= 159049 and INT_EDGE_VALUE <= 163591 else 
"01001000" when INT_EDGE_VALUE >= 163592 and INT_EDGE_VALUE <= 168199 else 
"01001001" when INT_EDGE_VALUE >= 168200 and INT_EDGE_VALUE <= 172871 else 
"01001010" when INT_EDGE_VALUE >= 172872 and INT_EDGE_VALUE <= 177608 else 
"01001011" when INT_EDGE_VALUE >= 177609 and INT_EDGE_VALUE <= 182407 else 
"01001100" when INT_EDGE_VALUE >= 182408 and INT_EDGE_VALUE <= 187271 else 
"01001101" when INT_EDGE_VALUE >= 187272 and INT_EDGE_VALUE <= 192199 else 
"01001110" when INT_EDGE_VALUE >= 192200 and INT_EDGE_VALUE <= 197191 else 
"01001111" when INT_EDGE_VALUE >= 197192 and INT_EDGE_VALUE <= 202247 else 
"01010000" when INT_EDGE_VALUE >= 202248 and INT_EDGE_VALUE <= 207367 else 
"01010001" when INT_EDGE_VALUE >= 207368 and INT_EDGE_VALUE <= 212551 else 
"01010010" when INT_EDGE_VALUE >= 212552 and INT_EDGE_VALUE <= 217799 else 
"01010011" when INT_EDGE_VALUE >= 217800 and INT_EDGE_VALUE <= 223111 else 
"01010100" when INT_EDGE_VALUE >= 223112 and INT_EDGE_VALUE <= 228487 else 
"01010101" when INT_EDGE_VALUE >= 228488 and INT_EDGE_VALUE <= 233927 else 
"01010110" when INT_EDGE_VALUE >= 233928 and INT_EDGE_VALUE <= 239432 else 
"01010111" when INT_EDGE_VALUE >= 239433 and INT_EDGE_VALUE <= 244999 else 
"01011000" when INT_EDGE_VALUE >= 245000 and INT_EDGE_VALUE <= 250631 else 
"01011001" when INT_EDGE_VALUE >= 250632 and INT_EDGE_VALUE <= 256327 else 
"01011010" when INT_EDGE_VALUE >= 256328 and INT_EDGE_VALUE <= 262088 else 
"01011011" when INT_EDGE_VALUE >= 262089 and INT_EDGE_VALUE <= 267912 else 
"01011100" when INT_EDGE_VALUE >= 267913 and INT_EDGE_VALUE <= 273799 else 
"01011101" when INT_EDGE_VALUE >= 273800 and INT_EDGE_VALUE <= 279751 else 
"01011110" when INT_EDGE_VALUE >= 279752 and INT_EDGE_VALUE <= 285768 else 
"01011111" when INT_EDGE_VALUE >= 285769 and INT_EDGE_VALUE <= 291847 else 
"01100000" when INT_EDGE_VALUE >= 291848 and INT_EDGE_VALUE <= 297991 else 
"01100001" when INT_EDGE_VALUE >= 297992 and INT_EDGE_VALUE <= 304199 else 
"01100010" when INT_EDGE_VALUE >= 304200 and INT_EDGE_VALUE <= 310472 else 
"01100011" when INT_EDGE_VALUE >= 310473 and INT_EDGE_VALUE <= 316807 else 
"01100100" when INT_EDGE_VALUE >= 316808 and INT_EDGE_VALUE <= 323207 else 
"01100101" when INT_EDGE_VALUE >= 323208 and INT_EDGE_VALUE <= 329671 else 
"01100110" when INT_EDGE_VALUE >= 329672 and INT_EDGE_VALUE <= 336199 else 
"01100111" when INT_EDGE_VALUE >= 336200 and INT_EDGE_VALUE <= 342792 else 
"01101000" when INT_EDGE_VALUE >= 342793 and INT_EDGE_VALUE <= 349447 else 
"01101001" when INT_EDGE_VALUE >= 349448 and INT_EDGE_VALUE <= 356167 else 
"01101010" when INT_EDGE_VALUE >= 356168 and INT_EDGE_VALUE <= 362952 else 
"01101011" when INT_EDGE_VALUE >= 362953 and INT_EDGE_VALUE <= 369799 else 
"01101100" when INT_EDGE_VALUE >= 369800 and INT_EDGE_VALUE <= 376712 else 
"01101101" when INT_EDGE_VALUE >= 376713 and INT_EDGE_VALUE <= 383687 else 
"01101110" when INT_EDGE_VALUE >= 383688 and INT_EDGE_VALUE <= 390727 else 
"01101111" when INT_EDGE_VALUE >= 390728 and INT_EDGE_VALUE <= 397832 else 
"01110000" when INT_EDGE_VALUE >= 397833 and INT_EDGE_VALUE <= 404999 else 
"01110001" when INT_EDGE_VALUE >= 405000 and INT_EDGE_VALUE <= 412231 else 
"01110010" when INT_EDGE_VALUE >= 412232 and INT_EDGE_VALUE <= 419528 else 
"01110011" when INT_EDGE_VALUE >= 419529 and INT_EDGE_VALUE <= 426887 else 
"01110100" when INT_EDGE_VALUE >= 426888 and INT_EDGE_VALUE <= 434311 else 
"01110101" when INT_EDGE_VALUE >= 434312 and INT_EDGE_VALUE <= 441799 else 
"01110110" when INT_EDGE_VALUE >= 441800 and INT_EDGE_VALUE <= 449352 else 
"01110111" when INT_EDGE_VALUE >= 449353 and INT_EDGE_VALUE <= 456967 else 
"01111000" when INT_EDGE_VALUE >= 456968 and INT_EDGE_VALUE <= 464647 else 
"01111001" when INT_EDGE_VALUE >= 464648 and INT_EDGE_VALUE <= 472391 else 
"01111010" when INT_EDGE_VALUE >= 472392 and INT_EDGE_VALUE <= 480199 else 
"01111011" when INT_EDGE_VALUE >= 480200 and INT_EDGE_VALUE <= 488072 else 
"01111100" when INT_EDGE_VALUE >= 488073 and INT_EDGE_VALUE <= 496007 else 
"01111101" when INT_EDGE_VALUE >= 496008 and INT_EDGE_VALUE <= 504007 else 
"01111110" when INT_EDGE_VALUE >= 504008 and INT_EDGE_VALUE <= 512072 else 
"01111111" when INT_EDGE_VALUE >= 512073 and INT_EDGE_VALUE <= 520199 else 
"10000000" when INT_EDGE_VALUE >= 520200 and INT_EDGE_VALUE <= 528391 else 
"10000001" when INT_EDGE_VALUE >= 528392 and INT_EDGE_VALUE <= 536647 else 
"10000010" when INT_EDGE_VALUE >= 536648 and INT_EDGE_VALUE <= 544967 else 
"10000011" when INT_EDGE_VALUE >= 544968 and INT_EDGE_VALUE <= 553351 else 
"10000100" when INT_EDGE_VALUE >= 553352 and INT_EDGE_VALUE <= 561799 else 
"10000101" when INT_EDGE_VALUE >= 561800 and INT_EDGE_VALUE <= 570312 else 
"10000110" when INT_EDGE_VALUE >= 570313 and INT_EDGE_VALUE <= 578887 else 
"10000111" when INT_EDGE_VALUE >= 578888 and INT_EDGE_VALUE <= 587527 else 
"10001000" when INT_EDGE_VALUE >= 587528 and INT_EDGE_VALUE <= 596231 else 
"10001001" when INT_EDGE_VALUE >= 596232 and INT_EDGE_VALUE <= 604999 else 
"10001010" when INT_EDGE_VALUE >= 605000 and INT_EDGE_VALUE <= 613831 else 
"10001011" when INT_EDGE_VALUE >= 613832 and INT_EDGE_VALUE <= 622728 else 
"10001100" when INT_EDGE_VALUE >= 622729 and INT_EDGE_VALUE <= 631687 else 
"10001101" when INT_EDGE_VALUE >= 631688 and INT_EDGE_VALUE <= 640712 else 
"10001110" when INT_EDGE_VALUE >= 640713 and INT_EDGE_VALUE <= 649799 else 
"10001111" when INT_EDGE_VALUE >= 649800 and INT_EDGE_VALUE <= 658951 else 
"10010000" when INT_EDGE_VALUE >= 658952 and INT_EDGE_VALUE <= 668167 else 
"10010001" when INT_EDGE_VALUE >= 668168 and INT_EDGE_VALUE <= 677447 else 
"10010010" when INT_EDGE_VALUE >= 677448 and INT_EDGE_VALUE <= 686791 else 
"10010011" when INT_EDGE_VALUE >= 686792 and INT_EDGE_VALUE <= 696199 else 
"10010100" when INT_EDGE_VALUE >= 696200 and INT_EDGE_VALUE <= 705672 else 
"10010101" when INT_EDGE_VALUE >= 705673 and INT_EDGE_VALUE <= 715207 else 
"10010110" when INT_EDGE_VALUE >= 715208 and INT_EDGE_VALUE <= 724807 else 
"10010111" when INT_EDGE_VALUE >= 724808 and INT_EDGE_VALUE <= 734471 else 
"10011000" when INT_EDGE_VALUE >= 734472 and INT_EDGE_VALUE <= 744199 else 
"10011001" when INT_EDGE_VALUE >= 744200 and INT_EDGE_VALUE <= 753991 else 
"10011010" when INT_EDGE_VALUE >= 753992 and INT_EDGE_VALUE <= 763847 else 
"10011011" when INT_EDGE_VALUE >= 763848 and INT_EDGE_VALUE <= 773767 else 
"10011100" when INT_EDGE_VALUE >= 773768 and INT_EDGE_VALUE <= 783752 else 
"10011101" when INT_EDGE_VALUE >= 783753 and INT_EDGE_VALUE <= 793799 else 
"10011110" when INT_EDGE_VALUE >= 793800 and INT_EDGE_VALUE <= 803912 else 
"10011111" when INT_EDGE_VALUE >= 803913 and INT_EDGE_VALUE <= 814087 else 
"10100000" when INT_EDGE_VALUE >= 814088 and INT_EDGE_VALUE <= 824327 else 
"10100001" when INT_EDGE_VALUE >= 824328 and INT_EDGE_VALUE <= 834631 else 
"10100010" when INT_EDGE_VALUE >= 834632 and INT_EDGE_VALUE <= 844999 else 
"10100011" when INT_EDGE_VALUE >= 845000 and INT_EDGE_VALUE <= 855432 else 
"10100100" when INT_EDGE_VALUE >= 855433 and INT_EDGE_VALUE <= 865927 else 
"10100101" when INT_EDGE_VALUE >= 865928 and INT_EDGE_VALUE <= 876488 else 
"10100110" when INT_EDGE_VALUE >= 876489 and INT_EDGE_VALUE <= 887111 else 
"10100111" when INT_EDGE_VALUE >= 887112 and INT_EDGE_VALUE <= 897799 else 
"10101000" when INT_EDGE_VALUE >= 897800 and INT_EDGE_VALUE <= 908551 else 
"10101001" when INT_EDGE_VALUE >= 908552 and INT_EDGE_VALUE <= 919367 else 
"10101010" when INT_EDGE_VALUE >= 919368 and INT_EDGE_VALUE <= 930247 else 
"10101011" when INT_EDGE_VALUE >= 930248 and INT_EDGE_VALUE <= 941192 else 
"10101100" when INT_EDGE_VALUE >= 941193 and INT_EDGE_VALUE <= 952199 else 
"10101101" when INT_EDGE_VALUE >= 952200 and INT_EDGE_VALUE <= 963272 else 
"10101110" when INT_EDGE_VALUE >= 963273 and INT_EDGE_VALUE <= 974407 else 
"10101111" when INT_EDGE_VALUE >= 974408 and INT_EDGE_VALUE <= 985608 else 
"10110000" when INT_EDGE_VALUE >= 985609 and INT_EDGE_VALUE <= 996871 else 
"10110001" when INT_EDGE_VALUE >= 996872 and INT_EDGE_VALUE <= 1008199 else 
"10110010" when INT_EDGE_VALUE >= 1008200 and INT_EDGE_VALUE <= 1019591 else 
"10110011" when INT_EDGE_VALUE >= 1019592 and INT_EDGE_VALUE <= 1031048 else 
"10110100" when INT_EDGE_VALUE >= 1031049 and INT_EDGE_VALUE <= 1042568 else 
"10110101" when INT_EDGE_VALUE >= 1042569 and INT_EDGE_VALUE <= 1054151 else 
"10110110" when INT_EDGE_VALUE >= 1054152 and INT_EDGE_VALUE <= 1065800 else 
"10110111" when INT_EDGE_VALUE >= 1065801 and INT_EDGE_VALUE <= 1077511 else 
"10111000" when INT_EDGE_VALUE >= 1077512 and INT_EDGE_VALUE <= 1089287 else 
"10111001" when INT_EDGE_VALUE >= 1089288 and INT_EDGE_VALUE <= 1101127 else 
"10111010" when INT_EDGE_VALUE >= 1101128 and INT_EDGE_VALUE <= 1113031 else 
"10111011" when INT_EDGE_VALUE >= 1113032 and INT_EDGE_VALUE <= 1125000 else 
"10111100" when INT_EDGE_VALUE >= 1125001 and INT_EDGE_VALUE <= 1137032 else 
"10111101" when INT_EDGE_VALUE >= 1137033 and INT_EDGE_VALUE <= 1149127 else 
"10111110" when INT_EDGE_VALUE >= 1149128 and INT_EDGE_VALUE <= 1161287 else 
"10111111" when INT_EDGE_VALUE >= 1161288 and INT_EDGE_VALUE <= 1173511 else 
"11000000" when INT_EDGE_VALUE >= 1173512 and INT_EDGE_VALUE <= 1185800 else 
"11000001" when INT_EDGE_VALUE >= 1185801 and INT_EDGE_VALUE <= 1198151 else 
"11000010" when INT_EDGE_VALUE >= 1198152 and INT_EDGE_VALUE <= 1210567 else 
"11000011" when INT_EDGE_VALUE >= 1210568 and INT_EDGE_VALUE <= 1223047 else 
"11000100" when INT_EDGE_VALUE >= 1223048 and INT_EDGE_VALUE <= 1235591 else 
"11000101" when INT_EDGE_VALUE >= 1235592 and INT_EDGE_VALUE <= 1248200 else 
"11000110" when INT_EDGE_VALUE >= 1248201 and INT_EDGE_VALUE <= 1260872 else 
"11000111" when INT_EDGE_VALUE >= 1260873 and INT_EDGE_VALUE <= 1273607 else 
"11001000" when INT_EDGE_VALUE >= 1273608 and INT_EDGE_VALUE <= 1286407 else 
"11001001" when INT_EDGE_VALUE >= 1286408 and INT_EDGE_VALUE <= 1299271 else 
"11001010" when INT_EDGE_VALUE >= 1299272 and INT_EDGE_VALUE <= 1312199 else 
"11001011" when INT_EDGE_VALUE >= 1312200 and INT_EDGE_VALUE <= 1325192 else 
"11001100" when INT_EDGE_VALUE >= 1325193 and INT_EDGE_VALUE <= 1338247 else 
"11001101" when INT_EDGE_VALUE >= 1338248 and INT_EDGE_VALUE <= 1351367 else 
"11001110" when INT_EDGE_VALUE >= 1351368 and INT_EDGE_VALUE <= 1364551 else 
"11001111" when INT_EDGE_VALUE >= 1364552 and INT_EDGE_VALUE <= 1377800 else 
"11010000" when INT_EDGE_VALUE >= 1377801 and INT_EDGE_VALUE <= 1391111 else 
"11010001" when INT_EDGE_VALUE >= 1391112 and INT_EDGE_VALUE <= 1404487 else 
"11010010" when INT_EDGE_VALUE >= 1404488 and INT_EDGE_VALUE <= 1417927 else 
"11010011" when INT_EDGE_VALUE >= 1417928 and INT_EDGE_VALUE <= 1431431 else 
"11010100" when INT_EDGE_VALUE >= 1431432 and INT_EDGE_VALUE <= 1445000 else 
"11010101" when INT_EDGE_VALUE >= 1445001 and INT_EDGE_VALUE <= 1458632 else 
"11010110" when INT_EDGE_VALUE >= 1458633 and INT_EDGE_VALUE <= 1472327 else 
"11010111" when INT_EDGE_VALUE >= 1472328 and INT_EDGE_VALUE <= 1486087 else 
"11011000" when INT_EDGE_VALUE >= 1486088 and INT_EDGE_VALUE <= 1499911 else 
"11011001" when INT_EDGE_VALUE >= 1499912 and INT_EDGE_VALUE <= 1513799 else 
"11011010" when INT_EDGE_VALUE >= 1513800 and INT_EDGE_VALUE <= 1527751 else 
"11011011" when INT_EDGE_VALUE >= 1527752 and INT_EDGE_VALUE <= 1541768 else 
"11011100" when INT_EDGE_VALUE >= 1541769 and INT_EDGE_VALUE <= 1555847 else 
"11011101" when INT_EDGE_VALUE >= 1555848 and INT_EDGE_VALUE <= 1569992 else 
"11011110" when INT_EDGE_VALUE >= 1569993 and INT_EDGE_VALUE <= 1584200 else 
"11011111" when INT_EDGE_VALUE >= 1584201 and INT_EDGE_VALUE <= 1598471 else 
"11100000" when INT_EDGE_VALUE >= 1598472 and INT_EDGE_VALUE <= 1612807 else 
"11100001" when INT_EDGE_VALUE >= 1612808 and INT_EDGE_VALUE <= 1627207 else 
"11100010" when INT_EDGE_VALUE >= 1627208 and INT_EDGE_VALUE <= 1641672 else 
"11100011" when INT_EDGE_VALUE >= 1641673 and INT_EDGE_VALUE <= 1656200 else 
"11100100" when INT_EDGE_VALUE >= 1656201 and INT_EDGE_VALUE <= 1670792 else 
"11100101" when INT_EDGE_VALUE >= 1670793 and INT_EDGE_VALUE <= 1685447 else 
"11100110" when INT_EDGE_VALUE >= 1685448 and INT_EDGE_VALUE <= 1700167 else 
"11100111" when INT_EDGE_VALUE >= 1700168 and INT_EDGE_VALUE <= 1714952 else 
"11101000" when INT_EDGE_VALUE >= 1714953 and INT_EDGE_VALUE <= 1729800 else 
"11101001" when INT_EDGE_VALUE >= 1729801 and INT_EDGE_VALUE <= 1744711 else 
"11101010" when INT_EDGE_VALUE >= 1744712 and INT_EDGE_VALUE <= 1759687 else 
"11101011" when INT_EDGE_VALUE >= 1759688 and INT_EDGE_VALUE <= 1774727 else 
"11101100" when INT_EDGE_VALUE >= 1774728 and INT_EDGE_VALUE <= 1789832 else 
"11101101" when INT_EDGE_VALUE >= 1789833 and INT_EDGE_VALUE <= 1805000 else 
"11101110" when INT_EDGE_VALUE >= 1805001 and INT_EDGE_VALUE <= 1820231 else 
"11101111" when INT_EDGE_VALUE >= 1820232 and INT_EDGE_VALUE <= 1835527 else 
"11110000" when INT_EDGE_VALUE >= 1835528 and INT_EDGE_VALUE <= 1850887 else 
"11110001" when INT_EDGE_VALUE >= 1850888 and INT_EDGE_VALUE <= 1866312 else 
"11110010" when INT_EDGE_VALUE >= 1866313 and INT_EDGE_VALUE <= 1881799 else 
"11110011" when INT_EDGE_VALUE >= 1881800 and INT_EDGE_VALUE <= 1897352 else 
"11110100" when INT_EDGE_VALUE >= 1897353 and INT_EDGE_VALUE <= 1912967 else 
"11110101" when INT_EDGE_VALUE >= 1912968 and INT_EDGE_VALUE <= 1928647 else 
"11110110" when INT_EDGE_VALUE >= 1928648 and INT_EDGE_VALUE <= 1944392 else 
"11110111" when INT_EDGE_VALUE >= 1944393 and INT_EDGE_VALUE <= 1960200 else 
"11111000" when INT_EDGE_VALUE >= 1960201 and INT_EDGE_VALUE <= 1976071 else 
"11111001" when INT_EDGE_VALUE >= 1976072 and INT_EDGE_VALUE <= 1992007 else 
"11111010" when INT_EDGE_VALUE >= 1992008 and INT_EDGE_VALUE <= 2008007 else 
"11111011" when INT_EDGE_VALUE >= 2008008 and INT_EDGE_VALUE <= 2024072 else 
"11111100" when INT_EDGE_VALUE >= 2024073 and INT_EDGE_VALUE <= 2040200 else 
"11111101" when INT_EDGE_VALUE >= 2040201 and INT_EDGE_VALUE <= 2056392 else 
"11111110" when INT_EDGE_VALUE >= 2056393 and INT_EDGE_VALUE <= 2072647 else 
"11111111" when INT_EDGE_VALUE >= 2072648; 

end architecture;